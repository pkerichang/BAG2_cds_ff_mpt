/tools/projects/jdhan/BAG/BAG2_cds_ff_mpt/pvs_run/netlist