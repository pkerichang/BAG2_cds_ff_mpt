** Layout Netlist, pvs precompare
** 

.subckt sar_wsamp ADCOUT<0> ADCOUT<1> ADCOUT<2> ADCOUT<3> ADCOUT<4> ADCOUT<5> ADCOUT<6> ADCOUT<7> ADCOUT<8> CKDSEL0<0> CKDSEL0<1> CKDSEL1<0> CKDSEL1<1> CLK CLKO CLKPRB_SAMP DONE EXTSEL_CLK ICLK INM 
+ INP OSM OSP PHI0 SAMPM SAMPP SAOM SAOP SARCLK SARCLKB SB<0> SB<1> SB<2> SB<3> SB<4> SB<5> SB<6> SB<7> SB<8> UP 
+ VDDSAMP VDDSAR VOL<0> VOL<1> VOL<2> VOL<3> VOL<4> VOL<5> VOL<6> VOL<7> VOR<0> VOR<1> VOR<2> VOR<3> VOR<4> VOR<5> VOR<6> VOR<7> VREF<0> VREF<1> 
+ VREF<2> VSS ZM<0> ZM<1> ZM<2> ZM<3> ZM<4> ZM<5> ZM<6> ZM<7> ZM<8> ZMID<0> ZMID<1> ZMID<2> ZMID<3> ZMID<4> ZMID<5> ZMID<7> ZP<0> ZP<1> 
+ ZP<3> ZP<4> ZP<5> ZP<7> ZP<8> 
RX81/X76/X50/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X51/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X52/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X53/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X54/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X55/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X56/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X57/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X58/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X59/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X60/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X61/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X62/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X63/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X64/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X65/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X66/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X67/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X68/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X69/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X70/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X71/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X72/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X73/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X74/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X75/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X76/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X77/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X78/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X79/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X80/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X81/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X82/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X83/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X84/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X85/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X86/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X87/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X88/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X89/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X90/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X91/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X92/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X93/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X94/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X95/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X96/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X97/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X98/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X99/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X100/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X101/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X102/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X103/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X104/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X105/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X106/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X107/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X108/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X109/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X110/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X111/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X112/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X113/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X114/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X115/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X116/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X117/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X118/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X119/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X120/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X121/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X122/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X123/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X124/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X125/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X126/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X127/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X128/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X129/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X130/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X131/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X132/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X133/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X134/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X135/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X136/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X137/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X138/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X139/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X140/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X141/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X142/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X143/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X144/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X145/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X146/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X147/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X148/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X149/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X150/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X151/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X152/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X153/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X154/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X155/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X156/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X157/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X158/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X159/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X160/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X161/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X162/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X163/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X164/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X165/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X166/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X167/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X168/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X169/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X170/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X171/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X172/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X173/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X174/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X175/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X176/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X177/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X178/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X179/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X180/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X181/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X182/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X183/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X184/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X185/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X186/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X187/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X188/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X189/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X190/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X191/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X192/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X193/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X194/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X195/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X196/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X197/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X198/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X199/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X200/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X201/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X202/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X203/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X204/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X205/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X206/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X207/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X208/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X209/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X210/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X211/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X212/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X213/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X214/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X215/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X216/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X217/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X218/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X219/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X220/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X221/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X222/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X223/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X224/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X225/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X226/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X227/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X228/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X229/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X230/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X231/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X232/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X233/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X234/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X235/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X236/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X237/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X238/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X239/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X240/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X241/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X242/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X243/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X244/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X245/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X246/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X247/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X248/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X249/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X250/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X251/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X252/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X253/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X254/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X255/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X256/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X257/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X258/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X259/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X260/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X261/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X76/X262/R0 SAMPP SAMPP RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X50/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X51/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X52/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X53/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X54/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X55/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X56/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X57/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X58/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X59/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X60/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X61/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X62/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X63/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X64/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X65/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X66/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X67/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X68/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X69/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X70/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X71/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X72/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X73/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X74/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X75/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X76/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X77/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X78/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X79/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X80/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X81/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X82/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X83/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X84/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X85/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X86/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X87/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X88/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X89/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X90/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X91/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X92/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X93/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X94/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X95/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X96/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X97/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X98/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X99/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X100/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X101/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X102/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X103/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X104/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X105/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X106/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X107/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X108/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X109/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X110/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X111/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X112/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X113/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X114/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X115/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X116/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X117/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X118/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X119/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X120/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X121/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X122/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X123/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X124/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X125/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X126/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X127/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X128/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X129/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X130/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X131/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X132/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X133/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X134/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X135/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X136/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X137/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X138/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X139/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X140/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X141/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X142/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X143/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X144/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X145/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X146/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X147/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X148/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X149/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X150/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X151/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X152/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X153/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X154/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X155/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X156/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X157/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X158/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X159/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X160/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X161/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X162/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X163/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X164/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X165/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X166/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X167/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X168/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X169/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X170/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X171/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X172/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X173/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X174/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X175/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X176/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X177/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X178/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X179/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X180/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X181/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X182/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X183/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X184/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X185/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X186/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X187/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X188/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X189/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X190/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X191/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X192/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X193/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X194/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X195/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X196/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X197/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X198/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X199/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X200/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X201/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X202/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X203/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X204/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X205/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X206/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X207/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X208/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X209/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X210/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X211/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X212/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X213/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X214/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X215/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X216/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X217/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X218/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X219/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X220/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X221/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X222/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X223/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X224/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X225/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X226/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X227/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X228/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X229/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X230/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X231/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X232/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X233/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X234/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X235/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X236/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X237/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X238/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X239/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X240/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X241/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X242/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X243/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X244/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X245/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X246/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X247/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X248/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X249/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X250/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X251/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X252/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X253/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X254/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X255/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X256/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X257/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X258/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X259/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X260/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X261/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
RX81/X77/X262/R0 SAMPM SAMPM RESM4 L=3.2e-08 W=3.2e-08 m=1 R=0.0604 
MX81/X86/X817/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X817/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X818/X0/M0 SAOP X81/X86/321 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X818/X1/M0 VDDSAR X81/X86/321 SAOP VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X819/X0/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X819/X1/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X820/X0/M0 SAOP X81/X86/321 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X820/X1/M0 VDDSAR X81/X86/321 SAOP VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X821/X0/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X821/X1/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X822/X0/M0 SAOP X81/X86/321 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X822/X1/M0 VDDSAR X81/X86/321 SAOP VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X823/X0/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X823/X1/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X824/X0/M0 SAOP X81/X86/321 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X824/X1/M0 VDDSAR X81/X86/321 SAOP VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X825/X0/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X825/X1/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X826/X0/M0 SAOP X81/X86/321 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X826/X1/M0 VDDSAR X81/X86/321 SAOP VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X827/X0/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X827/X1/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X828/X0/M0 SAOP X81/X86/321 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X828/X1/M0 VDDSAR X81/X86/321 SAOP VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X829/X0/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X829/X1/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X830/X0/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X830/X1/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X831/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X831/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X832/X0/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X832/X1/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X833/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X833/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X834/X0/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X834/X1/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X835/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X835/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X836/X0/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X836/X1/M0 VDDSAR OSP VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X837/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X837/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X838/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X838/X1/M0 X81/X86/324 VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X839/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X839/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X840/X0/M0 X81/397 OSP X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X840/X1/M0 X81/X86/324 OSP X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X841/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X841/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X842/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X842/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X843/X0/M0 X81/397 SAMPP X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X843/X1/M0 X81/X86/324 SAMPP X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X844/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X844/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X845/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X845/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X846/X0/M0 X81/397 SAMPP X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X846/X1/M0 X81/X86/324 SAMPP X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X847/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X847/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X848/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X848/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X849/X0/M0 X81/397 SAMPP X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X849/X1/M0 X81/X86/324 SAMPP X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X850/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X850/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X851/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X851/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X852/X0/M0 X81/397 SAMPP X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X852/X1/M0 X81/X86/324 SAMPP X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X853/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X853/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X854/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X854/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X855/X0/M0 X81/397 SAMPP X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X855/X1/M0 X81/X86/324 SAMPP X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X856/X0/M0 X81/X86/321 X81/X86/322 X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X856/X1/M0 X81/397 X81/X86/322 X81/X86/321 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X857/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X857/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X858/X0/M0 X81/397 SAMPP X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X858/X1/M0 X81/X86/324 SAMPP X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X859/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X859/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X860/X0/M0 X81/398 SAMPM X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X860/X1/M0 X81/X86/324 SAMPM X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X861/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X861/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X862/X0/M0 X81/398 SAMPM X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X862/X1/M0 X81/X86/324 SAMPM X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X863/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X863/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X864/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X864/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X865/X0/M0 X81/398 SAMPM X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X865/X1/M0 X81/X86/324 SAMPM X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X866/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X866/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X867/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X867/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X868/X0/M0 X81/398 SAMPM X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X868/X1/M0 X81/X86/324 SAMPM X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X869/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X869/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X870/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X870/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X871/X0/M0 X81/398 SAMPM X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X871/X1/M0 X81/X86/324 SAMPM X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X872/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X872/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X873/X0/M0 X81/X86/324 SARCLKB VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X873/X1/M0 VDDSAR SARCLKB X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X874/X0/M0 X81/398 SAMPM X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X874/X1/M0 X81/X86/324 SAMPM X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X875/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X875/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X876/X0/M0 X81/398 OSM X81/X86/324 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X876/X1/M0 X81/X86/324 OSM X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X877/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X877/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X878/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X878/X1/M0 X81/X86/324 VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X879/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X879/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X880/X0/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X880/X1/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X881/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X881/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X882/X0/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X882/X1/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X883/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X883/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X884/X0/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X884/X1/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X885/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X885/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X886/X0/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X886/X1/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X887/X0/M0 X81/X86/322 X81/X86/321 X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X887/X1/M0 X81/398 X81/X86/321 X81/X86/322 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X888/X0/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X888/X1/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X889/X0/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X889/X1/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X890/X0/M0 SAOM X81/X86/322 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X890/X1/M0 VDDSAR X81/X86/322 SAOM VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X891/X0/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X891/X1/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X892/X0/M0 SAOM X81/X86/322 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X892/X1/M0 VDDSAR X81/X86/322 SAOM VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X893/X0/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X893/X1/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X894/X0/M0 SAOM X81/X86/322 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X894/X1/M0 VDDSAR X81/X86/322 SAOM VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X895/X0/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X895/X1/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X896/X0/M0 SAOM X81/X86/322 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X896/X1/M0 VDDSAR X81/X86/322 SAOM VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X897/X0/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X897/X1/M0 VDDSAR OSM VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X898/X0/M0 SAOM X81/X86/322 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X898/X1/M0 VDDSAR X81/X86/322 SAOM VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X899/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X899/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X900/X0/M0 SAOM X81/X86/322 VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X900/X1/M0 VDDSAR X81/X86/322 SAOM VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1053/X4/M0 SAOP X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1053/X5/M0 VSS X81/X86/321 SAOP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1054/X4/M0 SAOP X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1054/X5/M0 VSS X81/X86/321 SAOP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1055/X4/M0 SAOP X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1055/X5/M0 VSS X81/X86/321 SAOP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1056/X4/M0 SAOP X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1056/X5/M0 VSS X81/X86/321 SAOP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1057/X4/M0 SAOP X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1057/X5/M0 VSS X81/X86/321 SAOP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1058/X4/M0 SAOP X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1058/X5/M0 VSS X81/X86/321 SAOP VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1059/X4/M0 X81/X86/321 X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1059/X5/M0 VSS X81/X86/322 X81/X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1060/X4/M0 X81/X86/321 X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1060/X5/M0 VSS X81/X86/322 X81/X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1061/X4/M0 X81/X86/321 X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1061/X5/M0 VSS X81/X86/322 X81/X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1062/X4/M0 X81/X86/321 X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1062/X5/M0 VSS X81/X86/322 X81/X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1063/X4/M0 X81/X86/321 X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1063/X5/M0 VSS X81/X86/322 X81/X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1064/X4/M0 X81/X86/321 X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1064/X5/M0 VSS X81/X86/322 X81/X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1065/X4/M0 X81/X86/321 X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1065/X5/M0 VSS X81/X86/322 X81/X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1066/X4/M0 X81/X86/321 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1066/X5/M0 VSS SARCLKB X81/X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1067/X4/M0 X81/X86/321 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1067/X5/M0 VSS SARCLKB X81/X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1068/X4/M0 X81/X86/321 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1068/X5/M0 VSS SARCLKB X81/X86/321 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1069/X4/M0 X81/397 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1069/X5/M0 VSS SARCLKB X81/397 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1070/X4/M0 X81/397 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1070/X5/M0 VSS SARCLKB X81/397 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1071/X4/M0 X81/397 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1071/X5/M0 VSS SARCLKB X81/397 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1072/X4/M0 X81/398 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1072/X5/M0 VSS SARCLKB X81/398 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1073/X4/M0 X81/398 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1073/X5/M0 VSS SARCLKB X81/398 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1074/X4/M0 X81/398 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1074/X5/M0 VSS SARCLKB X81/398 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1075/X4/M0 X81/X86/322 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1075/X5/M0 VSS SARCLKB X81/X86/322 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1076/X4/M0 X81/X86/322 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1076/X5/M0 VSS SARCLKB X81/X86/322 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1077/X4/M0 X81/X86/322 SARCLKB VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1077/X5/M0 VSS SARCLKB X81/X86/322 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1078/X4/M0 X81/X86/322 X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1078/X5/M0 VSS X81/X86/321 X81/X86/322 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1079/X4/M0 X81/X86/322 X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1079/X5/M0 VSS X81/X86/321 X81/X86/322 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1080/X4/M0 X81/X86/322 X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1080/X5/M0 VSS X81/X86/321 X81/X86/322 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1081/X4/M0 X81/X86/322 X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1081/X5/M0 VSS X81/X86/321 X81/X86/322 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1082/X4/M0 X81/X86/322 X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1082/X5/M0 VSS X81/X86/321 X81/X86/322 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1083/X4/M0 X81/X86/322 X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1083/X5/M0 VSS X81/X86/321 X81/X86/322 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1084/X4/M0 X81/X86/322 X81/X86/321 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1084/X5/M0 VSS X81/X86/321 X81/X86/322 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1085/X4/M0 SAOM X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1085/X5/M0 VSS X81/X86/322 SAOM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1086/X4/M0 SAOM X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1086/X5/M0 VSS X81/X86/322 SAOM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1087/X4/M0 SAOM X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1087/X5/M0 VSS X81/X86/322 SAOM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1088/X4/M0 SAOM X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1088/X5/M0 VSS X81/X86/322 SAOM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1089/X4/M0 SAOM X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1089/X5/M0 VSS X81/X86/322 SAOM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1090/X4/M0 SAOM X81/X86/322 VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1090/X5/M0 VSS X81/X86/322 SAOM VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1093/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1093/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1094/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1094/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1095/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1095/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1096/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1096/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1097/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1097/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1098/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1098/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1099/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1099/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1100/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1100/X1/M0 X81/397 VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1101/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1101/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1102/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1102/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1103/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1103/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1104/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1104/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1105/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1105/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1106/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1106/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1107/X0/M0 VDDSAR VDDSAR X81/397 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1107/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1108/X0/M0 VDDSAR VDDSAR X81/398 VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1108/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1109/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1109/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1110/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1110/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1111/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1111/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1112/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1112/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1113/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1113/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1114/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1114/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1115/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1115/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1116/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1116/X1/M0 X81/398 VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1117/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1117/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1118/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1118/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1119/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1119/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1120/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1120/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1121/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1121/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1122/X0/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX81/X86/X1122/X1/M0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X51/X0/M0 X82/X838/7 ICLK VDDSAR X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X51/X1/M0 VDDSAR ICLK X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X52/X0/M0 X82/X838/7 ICLK VDDSAR X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X52/X1/M0 VDDSAR ICLK X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X53/X0/M0 X82/X838/7 ICLK VDDSAR X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X53/X1/M0 VDDSAR ICLK X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X54/X0/M0 X82/X838/7 ICLK VDDSAR X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X54/X1/M0 VDDSAR ICLK X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X55/X0/M0 PHI0 X82/90 X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X55/X1/M0 X82/X838/7 X82/90 PHI0 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X56/X0/M0 PHI0 X82/90 X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X56/X1/M0 X82/X838/7 X82/90 PHI0 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X57/X0/M0 PHI0 X82/90 X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X57/X1/M0 X82/X838/7 X82/90 PHI0 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X58/X0/M0 PHI0 X82/90 X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X58/X1/M0 X82/X838/7 X82/90 PHI0 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X59/X0/M0 PHI0 DONE X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X59/X1/M0 X82/X838/7 DONE PHI0 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X60/X0/M0 PHI0 DONE X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X60/X1/M0 X82/X838/7 DONE PHI0 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X61/X0/M0 PHI0 DONE X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X61/X1/M0 X82/X838/7 DONE PHI0 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X62/X0/M0 PHI0 DONE X82/X838/7 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X62/X1/M0 X82/X838/7 DONE PHI0 X82/X838/9 P1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X63/X4/M0 PHI0 ICLK VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X63/X5/M0 VSS ICLK PHI0 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X64/X4/M0 X82/X838/13 X82/90 PHI0 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X64/X5/M0 PHI0 X82/90 X82/X838/13 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X65/X4/M0 X82/X838/13 X82/90 PHI0 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X65/X5/M0 PHI0 X82/90 X82/X838/13 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X66/X4/M0 X82/X838/13 X82/90 PHI0 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X66/X5/M0 PHI0 X82/90 X82/X838/13 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X67/X4/M0 X82/X838/13 X82/90 PHI0 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X67/X5/M0 PHI0 X82/90 X82/X838/13 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X68/X4/M0 X82/X838/13 DONE VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X68/X5/M0 VSS DONE X82/X838/13 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X69/X4/M0 X82/X838/13 DONE VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X69/X5/M0 VSS DONE X82/X838/13 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X70/X4/M0 X82/X838/13 DONE VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X70/X5/M0 VSS DONE X82/X838/13 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X71/X4/M0 X82/X838/13 DONE VSS VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
MX82/X838/X71/X5/M0 VSS DONE X82/X838/13 VSS N1LVT L=1.8e-08 nf=1 nfin=4 m=1 
.ends


