* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                          *
*                                                       *
* Cell Name  : latch_2ck_2x                             *
* Netlisted  : Thu Jun  1 20:55:23 2017                 *
* PVS Version: 15.17-s604 Fri Jun 24 15:14:35 PDT 2016 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: _nmos4_fast_base_nf1                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt _nmos4_fast_base_nf1 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 4 2 1 n1lvt L=1.8e-08 nf=1 nfin=4 $X=68 $Y=226
.ends _nmos4_fast_base_nf1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos4_fast_center_nf2                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos4_fast_center_nf2 S0 G0 D0 S1 5
** N=5 EP=5 FDC=2
X4 5 S0 D0 G0 _nmos4_fast_base_nf1 $T=0 0 0 0 $X=-234 $Y=-32
X5 5 D0 S1 G0 _nmos4_fast_base_nf1 $T=172 0 0 0 $X=-62 $Y=-32
.ends nmos4_fast_center_nf2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: _pmos4_fast_base_nf1                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt _pmos4_fast_base_nf1 1 3 4 5
** N=5 EP=4 FDC=1
M0 4 5 3 1 p1lvt L=1.8e-08 nf=1 nfin=4 $X=68 $Y=226
.ends _pmos4_fast_base_nf1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos4_fast_center_nf2                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos4_fast_center_nf2 S0 G0 D0 S1 5
** N=6 EP=5 FDC=2
X4 5 S0 D0 G0 _pmos4_fast_base_nf1 $T=0 0 0 0 $X=-234 $Y=-32
X5 5 D0 S1 G0 _pmos4_fast_base_nf1 $T=172 0 0 0 $X=-62 $Y=-32
.ends pmos4_fast_center_nf2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: tinv_2x                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt tinv_2x 1 I VSS VDD ENB O EN 10
** N=21 EP=8 FDC=8
X15 VSS I 11 VSS 1 nmos4_fast_center_nf2 $T=172 0 0 0 $X=-62 $Y=-32
X16 11 EN O 11 1 nmos4_fast_center_nf2 $T=860 0 0 0 $X=626 $Y=-32
X22 VDD I 12 VDD 10 pmos4_fast_center_nf2 $T=172 1920 1 0 $X=-62 $Y=928
X23 12 ENB O 12 10 pmos4_fast_center_nf2 $T=860 1920 1 0 $X=626 $Y=928
.ends tinv_2x

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inv_2x                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inv_2x 1 O I VSS VDD 8
** N=13 EP=6 FDC=4
X15 1 VSS O I _nmos4_fast_base_nf1 $T=172 0 0 0 $X=-62 $Y=-32
X16 1 O VSS I _nmos4_fast_base_nf1 $T=344 0 0 0 $X=110 $Y=-32
X24 8 VDD O I _pmos4_fast_base_nf1 $T=172 1920 1 0 $X=-62 $Y=928
X25 8 O VDD I _pmos4_fast_base_nf1 $T=344 1920 1 0 $X=110 $Y=928
.ends inv_2x

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: tinv_small_1x                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt tinv_small_1x 1 O I ENB VSS VDD EN 12
** N=22 EP=8 FDC=4
X11 1 VSS 13 I _nmos4_fast_base_nf1 $T=172 0 0 0 $X=-62 $Y=-32
X12 1 13 O EN _nmos4_fast_base_nf1 $T=344 0 0 0 $X=110 $Y=-32
X22 12 VDD 16 I _pmos4_fast_base_nf1 $T=172 1920 1 0 $X=-62 $Y=928
X23 12 16 O ENB _pmos4_fast_base_nf1 $T=344 1920 1 0 $X=110 $Y=928
.ends tinv_small_1x

* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: latch_2ck_2x                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt latch_2ck_2x CLK CLKB I O VDD VSS
** N=15 EP=6 FDC=16
X9 5 I VSS VDD CLKB 2 CLK 11 tinv_2x $T=0 0 0 0 $X=-104 $Y=-144
X10 5 O 2 VSS VDD 11 inv_2x $T=2408 0 0 0 $X=2304 $Y=-144
X11 5 2 O CLK VSS VDD CLKB 11 tinv_small_1x $T=1376 0 0 0 $X=1272 $Y=-144
.ends latch_2ck_2x
