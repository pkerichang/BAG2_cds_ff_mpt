** Schematic Netlist, pvs precompare
** 

.subckt sar_wsamp ADCOUT<8> ADCOUT<7> ADCOUT<6> ADCOUT<5> ADCOUT<4> ADCOUT<3> ADCOUT<2> ADCOUT<1> ADCOUT<0> CKDSEL0<1> CKDSEL0<0> CKDSEL1<1> CKDSEL1<0> CLK CLKO CLKPRB_SAMP DONE EXTSEL_CLK ICLK INM 
+ INP OSM OSP PHI0 SAMPM SAMPP SAOM SAOP SARCLK SARCLKB SB<8> SB<7> SB<6> SB<5> SB<4> SB<3> SB<2> SB<1> SB<0> UP 
+ VDDSAMP VDDSAR VOL<7> VOL<6> VOL<5> VOL<4> VOL<3> VOL<2> VOL<1> VOL<0> VOR<7> VOR<6> VOR<5> VOR<4> VOR<3> VOR<2> VOR<1> VOR<0> VREF<2> VREF<1> 
+ VREF<0> VSS ZM<8> ZM<7> ZM<6> ZM<5> ZM<4> ZM<3> ZM<2> ZM<1> ZM<0> ZMID<8> ZMID<7> ZMID<6> ZMID<5> ZMID<4> ZMID<3> ZMID<2> ZMID<1> ZMID<0> 
+ ZP<8> ZP<7> ZP<6> ZP<5> ZP<4> ZP<3> ZP<2> ZP<1> ZP<0> 
MXISAR0/XIABE0/XIRET0/XICKBUF3/XIN0/MM0 CLKO XISAR0/XIABE0/XIRET0/net06 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIABE0/XIRET0/XICKBUF3/XIP0/MM0 CLKO XISAR0/XIABE0/XIRET0/net06 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIABE0/XIRET0/XICKBUF1/XIN0/MM0 XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/net2 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIABE0/XIRET0/XICKBUF1/XIP0/MM0 XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/net2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIABE0/XIRET0/XICKBUF0/XIN0/MM0 XISAR0/XIABE0/XIRET0/net2 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XICKBUF0/XIP0/MM0 XISAR0/XIABE0/XIRET0/net2 ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XICKBUF2/XIN0/MM0 XISAR0/XIABE0/XIRET0/net06 XISAR0/XIABE0/XIRET0/ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XICKBUF2/XIP0/MM0 XISAR0/XIABE0/XIRET0/net06 XISAR0/XIABE0/XIRET0/ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI7/XIINV2/XIN0/MM0 ADCOUT<7> XISAR0/XIABE0/XIRET0/XI7/net12 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI7/XIINV2/XIP0/MM0 ADCOUT<7> XISAR0/XIABE0/XIRET0/XI7/net12 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI7/XIINV0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI7/CLKB XISAR0/XIABE0/XIRET0/ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XIINV0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI7/CLKB XISAR0/XIABE0/XIRET0/ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XIINV1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI7/net12 XISAR0/XIABE0/XIRET0/XI7/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XIINV1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI7/net12 XISAR0/XIABE0/XIRET0/XI7/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI7/net13 XISAR0/XIABE0/XIRET0/XI7/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI7/net13 XISAR0/XIABE0/XIRET0/XI7/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI7/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI0/N0 XISAR0/XIABE0/RETI<7> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI0/N1 XISAR0/XIABE0/RETI<7> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI7/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI7/CLKB XISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI7/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI7/CLKB XISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI2/N0 XISAR0/XIABE0/XIRET0/XI7/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI2/N1 XISAR0/XIABE0/XIRET0/XI7/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI7/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI7/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XIINV2/XIN0/MM0 ADCOUT<6> XISAR0/XIABE0/XIRET0/XI6/net12 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI6/XIINV2/XIP0/MM0 ADCOUT<6> XISAR0/XIABE0/XIRET0/XI6/net12 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI6/XIINV0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI6/CLKB XISAR0/XIABE0/XIRET0/ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XIINV0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI6/CLKB XISAR0/XIABE0/XIRET0/ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XIINV1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI6/net12 XISAR0/XIABE0/XIRET0/XI6/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XIINV1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI6/net12 XISAR0/XIABE0/XIRET0/XI6/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI6/net13 XISAR0/XIABE0/XIRET0/XI6/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI6/net13 XISAR0/XIABE0/XIRET0/XI6/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI6/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI0/N0 XISAR0/XIABE0/RETI<6> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI0/N1 XISAR0/XIABE0/RETI<6> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI6/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI6/CLKB XISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI6/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI6/CLKB XISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI2/N0 XISAR0/XIABE0/XIRET0/XI6/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI2/N1 XISAR0/XIABE0/XIRET0/XI6/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI6/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI6/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XIINV2/XIN0/MM0 ADCOUT<4> XISAR0/XIABE0/XIRET0/XI4/net12 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI4/XIINV2/XIP0/MM0 ADCOUT<4> XISAR0/XIABE0/XIRET0/XI4/net12 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI4/XIINV0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI4/CLKB XISAR0/XIABE0/XIRET0/ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XIINV0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI4/CLKB XISAR0/XIABE0/XIRET0/ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XIINV1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI4/net12 XISAR0/XIABE0/XIRET0/XI4/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XIINV1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI4/net12 XISAR0/XIABE0/XIRET0/XI4/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI4/net13 XISAR0/XIABE0/XIRET0/XI4/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI4/net13 XISAR0/XIABE0/XIRET0/XI4/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI4/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI0/N0 XISAR0/XIABE0/RETI<4> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI0/N1 XISAR0/XIABE0/RETI<4> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI4/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI4/CLKB XISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI4/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI4/CLKB XISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI2/N0 XISAR0/XIABE0/XIRET0/XI4/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI2/N1 XISAR0/XIABE0/XIRET0/XI4/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI4/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI4/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XIINV2/XIN0/MM0 ADCOUT<8> XISAR0/XIABE0/XIRET0/XI8/net12 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI8/XIINV2/XIP0/MM0 ADCOUT<8> XISAR0/XIABE0/XIRET0/XI8/net12 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI8/XIINV0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI8/CLKB XISAR0/XIABE0/XIRET0/ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XIINV0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI8/CLKB XISAR0/XIABE0/XIRET0/ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XIINV1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI8/net12 XISAR0/XIABE0/XIRET0/XI8/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XIINV1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI8/net12 XISAR0/XIABE0/XIRET0/XI8/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI8/net13 XISAR0/XIABE0/XIRET0/XI8/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI8/net13 XISAR0/XIABE0/XIRET0/XI8/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI8/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI0/N0 XISAR0/XIABE0/RETI<8> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI0/N1 XISAR0/XIABE0/RETI<8> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI8/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI8/CLKB XISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI8/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI8/CLKB XISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI2/N0 XISAR0/XIABE0/XIRET0/XI8/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI2/N1 XISAR0/XIABE0/XIRET0/XI8/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI8/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI8/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XIINV2/XIN0/MM0 ADCOUT<0> XISAR0/XIABE0/XIRET0/XI0/net12 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI0/XIINV2/XIP0/MM0 ADCOUT<0> XISAR0/XIABE0/XIRET0/XI0/net12 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI0/XIINV0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI0/CLKB XISAR0/XIABE0/XIRET0/ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XIINV0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI0/CLKB XISAR0/XIABE0/XIRET0/ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XIINV1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI0/net12 XISAR0/XIABE0/XIRET0/XI0/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XIINV1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI0/net12 XISAR0/XIABE0/XIRET0/XI0/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI0/net13 XISAR0/XIABE0/XIRET0/XI0/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI0/net13 XISAR0/XIABE0/XIRET0/XI0/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI0/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI0/N0 XISAR0/XIABE0/RETI<0> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI0/N1 XISAR0/XIABE0/RETI<0> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI0/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI0/CLKB XISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI0/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI0/CLKB XISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI2/N0 XISAR0/XIABE0/XIRET0/XI0/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI2/N1 XISAR0/XIABE0/XIRET0/XI0/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI0/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI0/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XIINV2/XIN0/MM0 ADCOUT<1> XISAR0/XIABE0/XIRET0/XI1/net12 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI1/XIINV2/XIP0/MM0 ADCOUT<1> XISAR0/XIABE0/XIRET0/XI1/net12 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI1/XIINV0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI1/CLKB XISAR0/XIABE0/XIRET0/ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XIINV0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI1/CLKB XISAR0/XIABE0/XIRET0/ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XIINV1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI1/net12 XISAR0/XIABE0/XIRET0/XI1/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XIINV1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI1/net12 XISAR0/XIABE0/XIRET0/XI1/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI1/net13 XISAR0/XIABE0/XIRET0/XI1/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI1/net13 XISAR0/XIABE0/XIRET0/XI1/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI1/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI0/N0 XISAR0/XIABE0/RETI<1> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI0/N1 XISAR0/XIABE0/RETI<1> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI1/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI1/CLKB XISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI1/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI1/CLKB XISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI2/N0 XISAR0/XIABE0/XIRET0/XI1/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI2/N1 XISAR0/XIABE0/XIRET0/XI1/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI1/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI1/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XIINV2/XIN0/MM0 ADCOUT<5> XISAR0/XIABE0/XIRET0/XI5/net12 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI5/XIINV2/XIP0/MM0 ADCOUT<5> XISAR0/XIABE0/XIRET0/XI5/net12 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI5/XIINV0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI5/CLKB XISAR0/XIABE0/XIRET0/ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XIINV0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI5/CLKB XISAR0/XIABE0/XIRET0/ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XIINV1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI5/net12 XISAR0/XIABE0/XIRET0/XI5/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XIINV1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI5/net12 XISAR0/XIABE0/XIRET0/XI5/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI5/net13 XISAR0/XIABE0/XIRET0/XI5/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI5/net13 XISAR0/XIABE0/XIRET0/XI5/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI5/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI0/N0 XISAR0/XIABE0/RETI<5> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI0/N1 XISAR0/XIABE0/RETI<5> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI5/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI5/CLKB XISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI5/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI5/CLKB XISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI2/N0 XISAR0/XIABE0/XIRET0/XI5/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI2/N1 XISAR0/XIABE0/XIRET0/XI5/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI5/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI5/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XIINV2/XIN0/MM0 ADCOUT<3> XISAR0/XIABE0/XIRET0/XI3/net12 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI3/XIINV2/XIP0/MM0 ADCOUT<3> XISAR0/XIABE0/XIRET0/XI3/net12 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI3/XIINV0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI3/CLKB XISAR0/XIABE0/XIRET0/ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XIINV0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI3/CLKB XISAR0/XIABE0/XIRET0/ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XIINV1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI3/net12 XISAR0/XIABE0/XIRET0/XI3/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XIINV1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI3/net12 XISAR0/XIABE0/XIRET0/XI3/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI3/net13 XISAR0/XIABE0/XIRET0/XI3/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI3/net13 XISAR0/XIABE0/XIRET0/XI3/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI3/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI0/N0 XISAR0/XIABE0/RETI<3> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI0/N1 XISAR0/XIABE0/RETI<3> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI3/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI3/CLKB XISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI3/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI3/CLKB XISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI2/N0 XISAR0/XIABE0/XIRET0/XI3/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI2/N1 XISAR0/XIABE0/XIRET0/XI3/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI3/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI3/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XIINV2/XIN0/MM0 ADCOUT<2> XISAR0/XIABE0/XIRET0/XI2/net12 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI2/XIINV2/XIP0/MM0 ADCOUT<2> XISAR0/XIABE0/XIRET0/XI2/net12 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XIRET0/XI2/XIINV0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI2/CLKB XISAR0/XIABE0/XIRET0/ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XIINV0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI2/CLKB XISAR0/XIABE0/XIRET0/ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XIINV1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI2/net12 XISAR0/XIABE0/XIRET0/XI2/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XIINV1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI2/net12 XISAR0/XIABE0/XIRET0/XI2/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI2/net13 XISAR0/XIABE0/XIRET0/XI2/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI2/net13 XISAR0/XIABE0/XIRET0/XI2/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI2/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI0/N0 XISAR0/XIABE0/RETI<2> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI0/N1 XISAR0/XIABE0/RETI<2> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI2/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI2/CLKB XISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XIRET0/XI2/XILATCH0/MEM XISAR0/XIABE0/XIRET0/XI2/CLKB XISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI2/N0 XISAR0/XIABE0/XIRET0/XI2/net13 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI2/N1 XISAR0/XIABE0/XIRET0/XI2/net13 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XIRET0/XI2/XILATCH0/MEM XISAR0/XIABE0/XIRET0/ICLK XISAR0/XIABE0/XIRET0/XI2/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/TRIGB XISAR0/XIABE0/RST_DLY VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/TRIGB XISAR0/XIABE0/RST_DLY VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI0/net6 XISAR0/XIABE0/XISARFSM0/XI0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI0/XIP0/MM0 VDDSAR XISAR0/XIABE0/XISARFSM0/XI0/net5 XISAR0/XIABE0/XISARFSM0/XI0/net5 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI7/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI7/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI6/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI6/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI8/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/IRSTB ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI8/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/IRSTB ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI5/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<0>/XI5/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI5/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI5/N0 SB<0> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI5/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI5/N1 SB<0> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI5/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<0>/XI5/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<0>/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI2/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI2/N0 XISAR0/XIABE0/XISARFSM0/XI3<0>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI2/N1 XISAR0/XIABE0/XISARFSM0/XI3<0>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI2/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<0>/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI4/XIN0/MM0 SB<0> XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI4/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI4/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI4/N0 XISAR0/XIABE0/XISARFSM0/XI3<0>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI4/XIP1/MM0 SB<0> XISAR0/XIABE0/XISARFSM0/XI3<0>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI4/XIP0/MM0 SB<0> XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI1/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI1/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI1/N0 XISAR0/XIABE0/XISARFSM0/XI3<0>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI1/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<0>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI1/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI3/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<0>/XI3/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI3/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI3/N0 XISAR0/XIABE0/XISARFSM0/XI3<0>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI3/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI3/N1 XISAR0/XIABE0/XISARFSM0/XI3<0>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI3/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<0>/XI3/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<0>/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI0/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI0/N0 SB<1> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI0/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/XI0/N1 SB<1> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<0>/XI0/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<0>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<0>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<0>/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI7/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI7/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI6/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI6/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI8/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/IRSTB ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI8/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/IRSTB ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI5/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<1>/XI5/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI5/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI5/N0 SB<1> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI5/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI5/N1 SB<1> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI5/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<1>/XI5/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<1>/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI2/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI2/N0 XISAR0/XIABE0/XISARFSM0/XI3<1>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI2/N1 XISAR0/XIABE0/XISARFSM0/XI3<1>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI2/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<1>/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI4/XIN0/MM0 SB<1> XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI4/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI4/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI4/N0 XISAR0/XIABE0/XISARFSM0/XI3<1>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI4/XIP1/MM0 SB<1> XISAR0/XIABE0/XISARFSM0/XI3<1>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI4/XIP0/MM0 SB<1> XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI1/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI1/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI1/N0 XISAR0/XIABE0/XISARFSM0/XI3<1>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI1/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<1>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI1/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI3/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<1>/XI3/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI3/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI3/N0 XISAR0/XIABE0/XISARFSM0/XI3<1>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI3/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI3/N1 XISAR0/XIABE0/XISARFSM0/XI3<1>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI3/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<1>/XI3/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<1>/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI0/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI0/N0 SB<2> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI0/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/XI0/N1 SB<2> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<1>/XI0/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<1>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<1>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<1>/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI7/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI7/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI6/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI6/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI8/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/IRSTB ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI8/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/IRSTB ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI5/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<2>/XI5/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI5/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI5/N0 SB<2> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI5/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI5/N1 SB<2> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI5/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<2>/XI5/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<2>/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI2/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI2/N0 XISAR0/XIABE0/XISARFSM0/XI3<2>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI2/N1 XISAR0/XIABE0/XISARFSM0/XI3<2>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI2/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<2>/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI4/XIN0/MM0 SB<2> XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI4/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI4/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI4/N0 XISAR0/XIABE0/XISARFSM0/XI3<2>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI4/XIP1/MM0 SB<2> XISAR0/XIABE0/XISARFSM0/XI3<2>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI4/XIP0/MM0 SB<2> XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI1/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI1/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI1/N0 XISAR0/XIABE0/XISARFSM0/XI3<2>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI1/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<2>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI1/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI3/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<2>/XI3/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI3/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI3/N0 XISAR0/XIABE0/XISARFSM0/XI3<2>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI3/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI3/N1 XISAR0/XIABE0/XISARFSM0/XI3<2>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI3/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<2>/XI3/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<2>/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI0/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI0/N0 SB<3> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI0/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/XI0/N1 SB<3> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<2>/XI0/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<2>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<2>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<2>/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI7/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI7/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI6/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI6/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI8/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/IRSTB ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI8/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/IRSTB ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI5/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<3>/XI5/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI5/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI5/N0 SB<3> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI5/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI5/N1 SB<3> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI5/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<3>/XI5/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<3>/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI2/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI2/N0 XISAR0/XIABE0/XISARFSM0/XI3<3>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI2/N1 XISAR0/XIABE0/XISARFSM0/XI3<3>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI2/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<3>/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI4/XIN0/MM0 SB<3> XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI4/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI4/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI4/N0 XISAR0/XIABE0/XISARFSM0/XI3<3>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI4/XIP1/MM0 SB<3> XISAR0/XIABE0/XISARFSM0/XI3<3>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI4/XIP0/MM0 SB<3> XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI1/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI1/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI1/N0 XISAR0/XIABE0/XISARFSM0/XI3<3>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI1/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<3>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI1/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI3/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<3>/XI3/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI3/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI3/N0 XISAR0/XIABE0/XISARFSM0/XI3<3>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI3/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI3/N1 XISAR0/XIABE0/XISARFSM0/XI3<3>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI3/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<3>/XI3/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<3>/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI0/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI0/N0 SB<4> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI0/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/XI0/N1 SB<4> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<3>/XI0/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<3>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<3>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<3>/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI7/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI7/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI6/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI6/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI8/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/IRSTB ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI8/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/IRSTB ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI5/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<4>/XI5/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI5/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI5/N0 SB<4> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI5/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI5/N1 SB<4> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI5/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<4>/XI5/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<4>/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI2/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI2/N0 XISAR0/XIABE0/XISARFSM0/XI3<4>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI2/N1 XISAR0/XIABE0/XISARFSM0/XI3<4>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI2/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<4>/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI4/XIN0/MM0 SB<4> XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI4/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI4/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI4/N0 XISAR0/XIABE0/XISARFSM0/XI3<4>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI4/XIP1/MM0 SB<4> XISAR0/XIABE0/XISARFSM0/XI3<4>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI4/XIP0/MM0 SB<4> XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI1/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI1/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI1/N0 XISAR0/XIABE0/XISARFSM0/XI3<4>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI1/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<4>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI1/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI3/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<4>/XI3/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI3/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI3/N0 XISAR0/XIABE0/XISARFSM0/XI3<4>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI3/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI3/N1 XISAR0/XIABE0/XISARFSM0/XI3<4>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI3/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<4>/XI3/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<4>/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI0/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI0/N0 SB<5> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI0/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/XI0/N1 SB<5> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<4>/XI0/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<4>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<4>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<4>/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI7/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI7/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI6/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI6/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI8/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/IRSTB ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI8/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/IRSTB ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI5/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<5>/XI5/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI5/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI5/N0 SB<5> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI5/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI5/N1 SB<5> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI5/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<5>/XI5/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<5>/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI2/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI2/N0 XISAR0/XIABE0/XISARFSM0/XI3<5>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI2/N1 XISAR0/XIABE0/XISARFSM0/XI3<5>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI2/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<5>/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI4/XIN0/MM0 SB<5> XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI4/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI4/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI4/N0 XISAR0/XIABE0/XISARFSM0/XI3<5>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI4/XIP1/MM0 SB<5> XISAR0/XIABE0/XISARFSM0/XI3<5>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI4/XIP0/MM0 SB<5> XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI1/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI1/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI1/N0 XISAR0/XIABE0/XISARFSM0/XI3<5>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI1/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<5>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI1/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI3/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<5>/XI3/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI3/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI3/N0 XISAR0/XIABE0/XISARFSM0/XI3<5>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI3/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI3/N1 XISAR0/XIABE0/XISARFSM0/XI3<5>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI3/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<5>/XI3/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<5>/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI0/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI0/N0 SB<6> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI0/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/XI0/N1 SB<6> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<5>/XI0/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<5>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<5>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<5>/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI7/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI7/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI6/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI6/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI8/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/IRSTB ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI8/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/IRSTB ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI5/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<6>/XI5/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI5/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI5/N0 SB<6> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI5/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI5/N1 SB<6> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI5/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<6>/XI5/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<6>/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI2/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI2/N0 XISAR0/XIABE0/XISARFSM0/XI3<6>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI2/N1 XISAR0/XIABE0/XISARFSM0/XI3<6>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI2/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<6>/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI4/XIN0/MM0 SB<6> XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI4/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI4/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI4/N0 XISAR0/XIABE0/XISARFSM0/XI3<6>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI4/XIP1/MM0 SB<6> XISAR0/XIABE0/XISARFSM0/XI3<6>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI4/XIP0/MM0 SB<6> XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI1/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI1/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI1/N0 XISAR0/XIABE0/XISARFSM0/XI3<6>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI1/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<6>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI1/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI3/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<6>/XI3/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI3/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI3/N0 XISAR0/XIABE0/XISARFSM0/XI3<6>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI3/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI3/N1 XISAR0/XIABE0/XISARFSM0/XI3<6>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI3/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<6>/XI3/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<6>/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI0/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI0/N0 SB<7> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI0/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/XI0/N1 SB<7> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<6>/XI0/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<6>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<6>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<6>/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI7/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI7/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI6/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI6/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI8/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/IRSTB ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI8/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/IRSTB ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI5/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<7>/XI5/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI5/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI5/N0 SB<7> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI5/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI5/N1 SB<7> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI5/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<7>/XI5/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<7>/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI2/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI2/N0 XISAR0/XIABE0/XISARFSM0/XI3<7>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI2/N1 XISAR0/XIABE0/XISARFSM0/XI3<7>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI2/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<7>/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI4/XIN0/MM0 SB<7> XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI4/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI4/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI4/N0 XISAR0/XIABE0/XISARFSM0/XI3<7>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI4/XIP1/MM0 SB<7> XISAR0/XIABE0/XISARFSM0/XI3<7>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI4/XIP0/MM0 SB<7> XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI1/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI1/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI1/N0 XISAR0/XIABE0/XISARFSM0/XI3<7>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI1/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<7>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI1/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI3/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<7>/XI3/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI3/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI3/N0 XISAR0/XIABE0/XISARFSM0/XI3<7>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI3/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI3/N1 XISAR0/XIABE0/XISARFSM0/XI3<7>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI3/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<7>/XI3/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<7>/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI0/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI0/N0 SB<8> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI0/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/XI0/N1 SB<8> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<7>/XI0/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<7>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<7>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<7>/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI7/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI7/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI6/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI6/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI8/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/IRSTB ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI8/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/IRSTB ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI5/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<8>/XI5/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI5/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI5/N0 SB<8> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI5/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI5/N1 SB<8> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI5/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<8>/XI5/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<8>/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI2/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI2/N0 XISAR0/XIABE0/XISARFSM0/XI3<8>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI2/N1 XISAR0/XIABE0/XISARFSM0/XI3<8>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI2/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<8>/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI4/XIN0/MM0 SB<8> XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI4/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI4/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI4/N0 XISAR0/XIABE0/XISARFSM0/XI3<8>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI4/XIP1/MM0 SB<8> XISAR0/XIABE0/XISARFSM0/XI3<8>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI4/XIP0/MM0 SB<8> XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI1/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI1/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI1/N0 XISAR0/XIABE0/XISARFSM0/XI3<8>/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI1/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<8>/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI1/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/LATCH XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI3/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<8>/XI3/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI3/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI3/N0 XISAR0/XIABE0/XISARFSM0/XI3<8>/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI3/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI3/N1 XISAR0/XIABE0/XISARFSM0/XI3<8>/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI3/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM2 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<8>/XI3/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLKB XISAR0/XIABE0/XISARFSM0/XI3<8>/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI0/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI0/N0 XISAR0/XIABE0/XISARFSM0/TRIGB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI0/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/XI0/N1 XISAR0/XIABE0/XISARFSM0/TRIGB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI3<8>/XI0/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI3<8>/MEM1 XISAR0/XIABE0/XISARFSM0/XI3<8>/ICLK XISAR0/XIABE0/XISARFSM0/XI3<8>/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI7/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/ICLK XISAR0/XIABE0/XISARFSM0/XI1/ICLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI7/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/ICLK XISAR0/XIABE0/XISARFSM0/XI1/ICLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI6/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/ICLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI6/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/ICLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI8/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/IRSTB ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI8/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/IRSTB ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI5/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/MEM2 XISAR0/XIABE0/XISARFSM0/XI1/ICLKB XISAR0/XIABE0/XISARFSM0/XI1/XI5/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI1/XI5/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/XI5/N0 XISAR0/XIABE0/RST_DLY VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI1/XI5/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/XI5/N1 XISAR0/XIABE0/RST_DLY VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI1/XI5/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/MEM2 XISAR0/XIABE0/XISARFSM0/XI1/ICLK XISAR0/XIABE0/XISARFSM0/XI1/XI5/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI1/XI2/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/MEM1 XISAR0/XIABE0/XISARFSM0/XI1/ICLK XISAR0/XIABE0/XISARFSM0/XI1/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI1/XI2/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/XI2/N0 XISAR0/XIABE0/XISARFSM0/XI1/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI1/XI2/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/XI2/N1 XISAR0/XIABE0/XISARFSM0/XI1/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI1/XI2/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/MEM1 XISAR0/XIABE0/XISARFSM0/XI1/ICLKB XISAR0/XIABE0/XISARFSM0/XI1/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARFSM0/XI1/XI4/XIN0/MM0 XISAR0/XIABE0/RST_DLY XISAR0/XIABE0/XISARFSM0/XI1/MEM2 XISAR0/XIABE0/XISARFSM0/XI1/XI4/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI4/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/XI4/N0 XISAR0/XIABE0/XISARFSM0/XI1/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI4/XIP1/MM0 XISAR0/XIABE0/RST_DLY XISAR0/XIABE0/XISARFSM0/XI1/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI4/XIP0/MM0 XISAR0/XIABE0/RST_DLY XISAR0/XIABE0/XISARFSM0/XI1/MEM2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI1/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/LATCH XISAR0/XIABE0/XISARFSM0/XI1/MEM1 XISAR0/XIABE0/XISARFSM0/XI1/XI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI1/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/XI1/N0 XISAR0/XIABE0/XISARFSM0/XI1/IRSTB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI1/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/LATCH XISAR0/XIABE0/XISARFSM0/XI1/IRSTB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI1/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/LATCH XISAR0/XIABE0/XISARFSM0/XI1/MEM1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI3/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/MEM2 XISAR0/XIABE0/XISARFSM0/XI1/ICLK XISAR0/XIABE0/XISARFSM0/XI1/XI3/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI3/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/XI3/N0 XISAR0/XIABE0/XISARFSM0/XI1/LATCH VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI3/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/XI3/N1 XISAR0/XIABE0/XISARFSM0/XI1/LATCH VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI3/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/MEM2 XISAR0/XIABE0/XISARFSM0/XI1/ICLKB XISAR0/XIABE0/XISARFSM0/XI1/XI3/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI0/XIN0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/MEM1 XISAR0/XIABE0/XISARFSM0/XI1/ICLKB XISAR0/XIABE0/XISARFSM0/XI1/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI0/XIN1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/XI0/N0 VSS VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI0/XIP0/MM0 XISAR0/XIABE0/XISARFSM0/XI1/XI0/N1 VSS VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARFSM0/XI1/XI0/XIP1/MM0 XISAR0/XIABE0/XISARFSM0/XI1/MEM1 XISAR0/XIABE0/XISARFSM0/XI1/ICLK XISAR0/XIABE0/XISARFSM0/XI1/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIINV0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/S SB<1> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIINV0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/S SB<1> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIINV3/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIINV3/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIINV2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIINV2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XINR0/XIN0/MM0 ZMID<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XINR0/XIN1/MM0 ZMID<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XINR0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XINR0/net04 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XINR0/XIP0/MM0 ZMID<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNOB XISAR0/XIABE0/XISARLOGIC0/XISL1/XINR0/net04 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNOB SB<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNOB SAOM XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/N0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/N3 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNOB SB<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNOB SB<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/N2 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/N1 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPOB SB<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPOB SAOP XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/N0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/N3 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPOB SB<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPOB SB<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/N2 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/N1 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL1/XIOAI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/RETI<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/RETI<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL1/S XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI0/N0 ZP<1> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI0/N1 ZP<1> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/MEM SB<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/MEM SB<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI2/N0 XISAR0/XIABE0/RETI<1> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI2/N1 XISAR0/XIABE0/RETI<1> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL1/S XISAR0/XIABE0/XISARLOGIC0/XISL1/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIBUF0/XIN0/MM0 ZM<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIBUF0/XIP0/MM0 ZM<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIBUF1/XIN0/MM0 ZP<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL1/XIBUF1/XIP0/MM0 ZP<1> XISAR0/XIABE0/XISARLOGIC0/XISL1/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIINV0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/S SB<2> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIINV0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/S SB<2> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIINV3/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIINV3/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIINV2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIINV2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XINR0/XIN0/MM0 ZMID<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XINR0/XIN1/MM0 ZMID<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XINR0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XINR0/net04 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XINR0/XIP0/MM0 ZMID<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNOB XISAR0/XIABE0/XISARLOGIC0/XISL2/XINR0/net04 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNOB SB<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNOB SAOM XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/N0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/N3 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNOB SB<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNOB SB<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/N2 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/N1 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPOB SB<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPOB SAOP XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/N0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/N3 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPOB SB<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPOB SB<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/N2 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/N1 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL2/XIOAI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/RETI<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/RETI<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL2/S XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI0/N0 ZP<2> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI0/N1 ZP<2> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/MEM SB<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/MEM SB<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI2/N0 XISAR0/XIABE0/RETI<2> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI2/N1 XISAR0/XIABE0/RETI<2> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL2/S XISAR0/XIABE0/XISARLOGIC0/XISL2/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIBUF0/XIN0/MM0 ZM<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIBUF0/XIP0/MM0 ZM<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIBUF1/XIN0/MM0 ZP<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL2/XIBUF1/XIP0/MM0 ZP<2> XISAR0/XIABE0/XISARLOGIC0/XISL2/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIINV0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/S SB<3> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIINV0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/S SB<3> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIINV3/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIINV3/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIINV2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIINV2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XINR0/XIN0/MM0 ZMID<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XINR0/XIN1/MM0 ZMID<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XINR0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XINR0/net04 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XINR0/XIP0/MM0 ZMID<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNOB XISAR0/XIABE0/XISARLOGIC0/XISL3/XINR0/net04 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNOB SB<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNOB SAOM XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/N0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/N3 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNOB SB<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNOB SB<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/N2 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/N1 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPOB SB<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPOB SAOP XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/N0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/N3 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPOB SB<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPOB SB<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/N2 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/N1 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL3/XIOAI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/RETI<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/RETI<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL3/S XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI0/N0 ZP<3> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI0/N1 ZP<3> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/MEM SB<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/MEM SB<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI2/N0 XISAR0/XIABE0/RETI<3> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI2/N1 XISAR0/XIABE0/RETI<3> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL3/S XISAR0/XIABE0/XISARLOGIC0/XISL3/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIBUF0/XIN0/MM0 ZM<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIBUF0/XIP0/MM0 ZM<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIBUF1/XIN0/MM0 ZP<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL3/XIBUF1/XIP0/MM0 ZP<3> XISAR0/XIABE0/XISARLOGIC0/XISL3/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIINV0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/S SB<4> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIINV0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/S SB<4> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIINV3/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIINV3/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIINV2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIINV2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XINR0/XIN0/MM0 ZMID<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XINR0/XIN1/MM0 ZMID<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XINR0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XINR0/net04 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XINR0/XIP0/MM0 ZMID<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNOB XISAR0/XIABE0/XISARLOGIC0/XISL4/XINR0/net04 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNOB SB<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNOB SAOM XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/N0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/N3 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNOB SB<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNOB SB<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/N2 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/N1 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPOB SB<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPOB SAOP XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/N0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/N3 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPOB SB<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPOB SB<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/N2 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/N1 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL4/XIOAI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/RETI<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/RETI<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL4/S XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI0/N0 ZP<4> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI0/N1 ZP<4> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/MEM SB<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/MEM SB<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI2/N0 XISAR0/XIABE0/RETI<4> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI2/N1 XISAR0/XIABE0/RETI<4> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL4/S XISAR0/XIABE0/XISARLOGIC0/XISL4/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIBUF0/XIN0/MM0 ZM<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIBUF0/XIP0/MM0 ZM<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIBUF1/XIN0/MM0 ZP<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL4/XIBUF1/XIP0/MM0 ZP<4> XISAR0/XIABE0/XISARLOGIC0/XISL4/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIINV0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/S SB<5> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIINV0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/S SB<5> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIINV3/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIINV3/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIINV2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIINV2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XINR0/XIN0/MM0 ZMID<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XINR0/XIN1/MM0 ZMID<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XINR0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XINR0/net04 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XINR0/XIP0/MM0 ZMID<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNOB XISAR0/XIABE0/XISARLOGIC0/XISL5/XINR0/net04 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNOB SB<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNOB SAOM XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/N0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/N3 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNOB SB<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNOB SB<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/N2 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/N1 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPOB SB<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPOB SAOP XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/N0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/N3 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPOB SB<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPOB SB<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/N2 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/N1 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL5/XIOAI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/RETI<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/RETI<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL5/S XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI0/N0 ZP<5> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI0/N1 ZP<5> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/MEM SB<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/MEM SB<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI2/N0 XISAR0/XIABE0/RETI<5> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI2/N1 XISAR0/XIABE0/RETI<5> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL5/S XISAR0/XIABE0/XISARLOGIC0/XISL5/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIBUF0/XIN0/MM0 ZM<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIBUF0/XIP0/MM0 ZM<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIBUF1/XIN0/MM0 ZP<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL5/XIBUF1/XIP0/MM0 ZP<5> XISAR0/XIABE0/XISARLOGIC0/XISL5/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIINV0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/S SB<6> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIINV0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/S SB<6> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIINV3/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIINV3/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIINV2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIINV2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XINR0/XIN0/MM0 ZMID<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XINR0/XIN1/MM0 ZMID<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XINR0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XINR0/net04 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XINR0/XIP0/MM0 ZMID<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNOB XISAR0/XIABE0/XISARLOGIC0/XISL6/XINR0/net04 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNOB SB<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNOB SAOM XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/N0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/N3 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNOB SB<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNOB SB<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/N2 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/N1 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPOB SB<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPOB SAOP XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/N0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/N3 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPOB SB<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPOB SB<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/N2 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/N1 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL6/XIOAI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/RETI<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/RETI<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL6/S XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI0/N0 ZP<6> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI0/N1 ZP<6> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/MEM SB<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/MEM SB<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI2/N0 XISAR0/XIABE0/RETI<6> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI2/N1 XISAR0/XIABE0/RETI<6> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL6/S XISAR0/XIABE0/XISARLOGIC0/XISL6/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIBUF0/XIN0/MM0 ZM<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIBUF0/XIP0/MM0 ZM<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIBUF1/XIN0/MM0 ZP<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL6/XIBUF1/XIP0/MM0 ZP<6> XISAR0/XIABE0/XISARLOGIC0/XISL6/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIINV0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/S SB<7> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIINV0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/S SB<7> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIINV3/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIINV3/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIINV2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIINV2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XINR0/XIN0/MM0 ZMID<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XINR0/XIN1/MM0 ZMID<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XINR0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XINR0/net04 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XINR0/XIP0/MM0 ZMID<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNOB XISAR0/XIABE0/XISARLOGIC0/XISL7/XINR0/net04 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNOB SB<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNOB SAOM XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/N0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/N3 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNOB SB<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNOB SB<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/N2 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/N1 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPOB SB<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPOB SAOP XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/N0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/N3 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPOB SB<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPOB SB<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/N2 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/N1 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL7/XIOAI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/RETI<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/RETI<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL7/S XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI0/N0 ZP<7> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI0/N1 ZP<7> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/MEM SB<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/MEM SB<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI2/N0 XISAR0/XIABE0/RETI<7> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI2/N1 XISAR0/XIABE0/RETI<7> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL7/S XISAR0/XIABE0/XISARLOGIC0/XISL7/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIBUF0/XIN0/MM0 ZM<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIBUF0/XIP0/MM0 ZM<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIBUF1/XIN0/MM0 ZP<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL7/XIBUF1/XIP0/MM0 ZP<7> XISAR0/XIABE0/XISARLOGIC0/XISL7/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIINV0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/S SB<0> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIINV0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/S SB<0> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIINV3/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIINV3/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIINV2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIINV2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XINR0/XIN0/MM0 ZMID<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XINR0/XIN1/MM0 ZMID<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XINR0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XINR0/net04 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XINR0/XIP0/MM0 ZMID<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNOB XISAR0/XIABE0/XISARLOGIC0/XISL0/XINR0/net04 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNOB SB<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNOB SAOM XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/N0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/N3 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNOB SB<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNOB SB<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/N2 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/N1 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPOB SB<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPOB SAOP XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/N0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/N3 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPOB SB<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPOB SB<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/N2 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/N1 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL0/XIOAI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/RETI<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/RETI<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL0/S XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI0/N0 ZP<0> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI0/N1 ZP<0> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/MEM SB<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/MEM SB<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI2/N0 XISAR0/XIABE0/RETI<0> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI2/N1 XISAR0/XIABE0/RETI<0> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL0/S XISAR0/XIABE0/XISARLOGIC0/XISL0/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIBUF0/XIN0/MM0 ZM<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIBUF0/XIP0/MM0 ZM<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIBUF1/XIN0/MM0 ZP<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL0/XIBUF1/XIP0/MM0 ZP<0> XISAR0/XIABE0/XISARLOGIC0/XISL0/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIINV0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/S SB<8> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIINV0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/S SB<8> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIINV3/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIINV3/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNO XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIINV2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIINV2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPO XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XINR0/XIN0/MM0 ZMID<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XINR0/XIN1/MM0 ZMID<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPOB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XINR0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XINR0/net04 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPOB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XINR0/XIP0/MM0 ZMID<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNOB XISAR0/XIABE0/XISARLOGIC0/XISL8/XINR0/net04 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNOB SB<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNOB SAOM XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/N0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/N3 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNOB SB<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNOB SB<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/N2 SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/N1 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/XIN2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPOB SB<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/XIN3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/N0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPOB SAOP XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/N0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/XIP4/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/N3 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/XIP5/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPOB SB<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/N3 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/XIP3/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPOB SB<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/N2 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/XIP2/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/N2 SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/N1 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPOB ICLK XISAR0/XIABE0/XISARLOGIC0/XISL8/XIOAI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI1/XIN0/MM0 XISAR0/XIABE0/RETI<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/MEM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI1/XIP0/MM0 XISAR0/XIABE0/RETI<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/MEM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI0/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL8/S XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI0/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI0/N0 ZP<8> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI0/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI0/N1 ZP<8> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI0/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/MEM SB<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI2/XIN0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/MEM SB<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI2/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI2/XIN1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI2/N0 XISAR0/XIABE0/RETI<8> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI2/XIP0/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI2/N1 XISAR0/XIABE0/RETI<8> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI2/XIP1/MM0 XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/MEM XISAR0/XIABE0/XISARLOGIC0/XISL8/S XISAR0/XIABE0/XISARLOGIC0/XISL8/XILATCH0/XI2/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIBUF0/XIN0/MM0 ZM<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIBUF0/XIP0/MM0 ZM<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/LDPO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIBUF1/XIN0/MM0 ZP<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNO VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XISARLOGIC0/XISL8/XIBUF1/XIP0/MM0 ZP<8> XISAR0/XIABE0/XISARLOGIC0/XISL8/LDNO VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XICKGEN0/XIINV8/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/CLKB PHI0 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIABE0/XICKGEN0/XIINV8/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/CLKB PHI0 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIABE0/XICKGEN0/XIINV5/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/UPB UP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XICKGEN0/XIINV5/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/UPB UP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XICKGEN0/XIINV1/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/SELINV<1> CKDSEL0<1> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIINV1/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/SELINV<1> CKDSEL0<1> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIINV0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/SELINV<0> CKDSEL0<0> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIINV0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/SELINV<0> CKDSEL0<0> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIINV2/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/SELINV<2> CKDSEL1<0> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIINV2/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/SELINV<2> CKDSEL1<0> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIINV7/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/EXTSELB_CLK EXTSEL_CLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIINV7/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/EXTSELB_CLK EXTSEL_CLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIINV0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN1 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN0 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIINV0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN1 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN0 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XINR0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN0 ZMID<6> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XINR0/XIN1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN0 XISAR0/XIABE0/XICKGEN0/EXTSELB_CLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XINR0/XIP1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XINR0/net04 XISAR0/XIABE0/XICKGEN0/EXTSELB_CLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XINR0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN0 ZMID<6> XISAR0/XIABE0/XICKGEN0/XIDLY0/XINR0/net04 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XIINV0/XIN0/MM0 UP XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/net8 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XIINV0/XIP0/MM0 UP XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/net8 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV1/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN1 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV1/XIN1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV1/N0 XISAR0/XIABE0/XICKGEN0/XIDLY0/n2 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV1/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV1/N1 XISAR0/XIABE0/XICKGEN0/XIDLY0/n2 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV1/XIP1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV0/XIN1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV0/N0 XISAR0/XIABE0/XICKGEN0/XIDLY0/n0 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV0/N1 XISAR0/XIABE0/XICKGEN0/XIDLY0/n0 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV0/XIP1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/XIDLY0/EN1 XISAR0/XIABE0/XICKGEN0/XIDLY0/XIMUX0/XITINV0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIINVSEL0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/SELB XISAR0/XIABE0/XICKGEN0/SELINV<0> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIINVSEL0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/SELB XISAR0/XIABE0/XICKGEN0/SELINV<0> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIINVDB0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/CKD1 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/INT<1> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIINVDB0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/CKD1 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/INT<1> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIINVDA0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/INT<1> DONE VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIINVDA0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/INT<1> DONE VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XIINV0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/n0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/net8 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XIINV0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/n0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/net8 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV1/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/SELINV<0> XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV1/XIN1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV1/N0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/CKD1 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV1/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV1/N1 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/CKD1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV1/XIP1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/SELB XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/SELB XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV0/XIN1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV0/N0 DONE VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV0/N1 DONE VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV0/XIP1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/SELINV<0> XISAR0/XIABE0/XICKGEN0/XIDLY0/XI0/XIMUX0/XITINV0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIINVSEL0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/SELB XISAR0/XIABE0/XICKGEN0/SELINV<1> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIINVSEL0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/SELB XISAR0/XIABE0/XICKGEN0/SELINV<1> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIINVDB0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/CKD1 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/INT<1> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIINVDB0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/CKD1 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/INT<1> VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIINVDA0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/INT<1> XISAR0/XIABE0/XICKGEN0/XIDLY0/n0 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIINVDA0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/INT<1> XISAR0/XIABE0/XICKGEN0/XIDLY0/n0 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XIINV0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/n2 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/net8 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XIINV0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/n2 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/net8 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV1/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/SELINV<1> XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV1/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV1/XIN1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV1/N0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/CKD1 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV1/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV1/N1 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/CKD1 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV1/XIP1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/SELB XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV1/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV0/XIN0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/SELB XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV0/XIN1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV0/N0 XISAR0/XIABE0/XICKGEN0/XIDLY0/n0 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV0/N1 XISAR0/XIABE0/XICKGEN0/XIDLY0/n0 VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV0/XIP1/MM0 XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/net8 XISAR0/XIABE0/XICKGEN0/SELINV<1> XISAR0/XIABE0/XICKGEN0/XIDLY0/XI1/XIMUX0/XITINV0/N1 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=1 
MXISAR0/XIABE0/XICKGEN0/XIINV8C/XIN0/MM0 SARCLKB SARCLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=16 
MXISAR0/XIABE0/XICKGEN0/XIINV8C/XIP0/MM0 SARCLKB SARCLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=16 
MXISAR0/XIABE0/XICKGEN0/XIINV8B/XIN0/MM0 SARCLK XISAR0/XIABE0/XICKGEN0/CLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=16 
MXISAR0/XIABE0/XICKGEN0/XIINV8B/XIP0/MM0 SARCLK XISAR0/XIABE0/XICKGEN0/CLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=16 
MXISAR0/XIABE0/XICKGEN0/XIND0/XIN0/MM0 DONE SAOP XISAR0/XIABE0/XICKGEN0/XIND0/N0 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XICKGEN0/XIND0/XIN1/MM0 XISAR0/XIABE0/XICKGEN0/XIND0/N0 SAOM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XICKGEN0/XIND0/XIP1/MM0 DONE SAOM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XICKGEN0/XIND0/XIP0/MM0 DONE SAOP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIABE0/XICKGEN0/XICORE0/XIN2/MM0 XISAR0/XIABE0/XICKGEN0/XICORE0/net017 DONE VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIABE0/XICKGEN0/XICORE0/XIN0/MM0 PHI0 ICLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIABE0/XICKGEN0/XICORE0/XIN1/MM0 PHI0 XISAR0/XIABE0/XICKGEN0/UPB XISAR0/XIABE0/XICKGEN0/XICORE0/net017 VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIABE0/XICKGEN0/XICORE0/XIP2/MM0 PHI0 DONE XISAR0/XIABE0/XICKGEN0/XICORE0/net03 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIABE0/XICKGEN0/XICORE0/XIP0/MM0 XISAR0/XIABE0/XICKGEN0/XICORE0/net03 ICLK VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIABE0/XICKGEN0/XICORE0/XIP1/MM0 PHI0 XISAR0/XIABE0/XICKGEN0/UPB XISAR0/XIABE0/XICKGEN0/XICORE0/net03 VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XISA0/XIRGNNDM1/MM0 XISAR0/XIAFE0/XISA0/OP XISAR0/XIAFE0/XISA0/OM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XISA0/XIBUFN0/MM0 SAOP XISAR0/XIAFE0/XISA0/OM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISAR0/XIAFE0/XISA0/XIBUFN1/MM0 SAOM XISAR0/XIAFE0/XISA0/OP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISAR0/XIAFE0/XISA0/XIRST1/MM0 XISAR0/XIAFE0/INTP SARCLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISAR0/XIAFE0/XISA0/XIRST3/MM0 XISAR0/XIAFE0/XISA0/OP SARCLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISAR0/XIAFE0/XISA0/XIRST0/MM0 XISAR0/XIAFE0/INTM SARCLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISAR0/XIAFE0/XISA0/XIRST2/MM0 XISAR0/XIAFE0/XISA0/OM SARCLKB VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISAR0/XIAFE0/XISA0/XIRGNNDM0/MM0 XISAR0/XIAFE0/XISA0/OM XISAR0/XIAFE0/XISA0/OP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XISA0/XIRGNN0/MM0 XISAR0/XIAFE0/XISA0/OM XISAR0/XIAFE0/XISA0/OP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISAR0/XIAFE0/XISA0/XIRGNN1/MM0 XISAR0/XIAFE0/XISA0/OP XISAR0/XIAFE0/XISA0/OM VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISAR0/XIAFE0/XISA0/XIBUFP0/MM0 SAOP XISAR0/XIAFE0/XISA0/OM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISAR0/XIAFE0/XISA0/XIBUFP1/MM0 SAOM XISAR0/XIAFE0/XISA0/OP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISAR0/XIAFE0/XISA0/XIRGNPDM2/MM0 XISAR0/XIAFE0/INTP VDDSAR VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XISA0/XIRGNPDM1/MM0 XISAR0/XIAFE0/INTM VDDSAR VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XISA0/XIRGNPDM0/MM0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XISA0/XIRGNP1/MM0 XISAR0/XIAFE0/XISA0/OP XISAR0/XIAFE0/XISA0/OM XISAR0/XIAFE0/INTP VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=22 
MXISAR0/XIAFE0/XISA0/XIRGNP0/MM0 XISAR0/XIAFE0/XISA0/OM XISAR0/XIAFE0/XISA0/OP XISAR0/XIAFE0/INTM VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=22 
MXISAR0/XIAFE0/XISA0/XIOSM0/MM0 XISAR0/XIAFE0/INTP OSM XISAR0/XIAFE0/XISA0/TAIL VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XISA0/XIOSP0/MM0 XISAR0/XIAFE0/INTM OSP XISAR0/XIAFE0/XISA0/TAIL VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XISA0/XIOSPB0/MM0 VDDSAR OSP VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=20 
MXISAR0/XIAFE0/XISA0/XIOSMB0/MM0 VDDSAR OSM VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=20 
MXISAR0/XIAFE0/XISA0/XIINDM1/MM0 VDDSAR VDDSAR XISAR0/XIAFE0/XISA0/TAIL VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XISA0/XIINDM0/MM0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=6 
MXISAR0/XIAFE0/XISA0/XICKPDM0/MM0 VDDSAR VDDSAR VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=52 
MXISAR0/XIAFE0/XISA0/XICKP0/MM0 XISAR0/XIAFE0/XISA0/TAIL SARCLKB VDDSAR VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=24 
MXISAR0/XIAFE0/XISA0/XIINM0/MM0 XISAR0/XIAFE0/INTP SAMPM XISAR0/XIAFE0/XISA0/TAIL VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISAR0/XIAFE0/XISA0/XIINP0/MM0 XISAR0/XIAFE0/INTM SAMPP XISAR0/XIAFE0/XISA0/TAIL VDDSAR P1LVT m=1 l=1.8e-08 nfin=4 nf=12 
MXISAR0/XIAFE0/XICDRVM0/XICDRV3/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV3/XITIE0/net5 XISAR0/XIAFE0/XICDRVM0/XICDRV3/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV3/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV3/XITIE0/net6 XISAR0/XIAFE0/XICDRVM0/XICDRV3/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV3/XISW0/XIN1/MM0 VREF<2> ZP<4> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV3/XISW0/XIN0/MM0 VREF<2> ZP<4> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV3/XISW1/XIN1/MM0 VREF<1> ZMID<4> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV3/XISW1/XIN0/MM0 VREF<1> ZMID<4> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV3/XISW2/XIN1/MM0 VREF<0> ZM<4> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV3/XISW2/XIN0/MM0 VREF<0> ZM<4> VOR<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV0/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV0/XITIE0/net5 XISAR0/XIAFE0/XICDRVM0/XICDRV0/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV0/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV0/XITIE0/net6 XISAR0/XIAFE0/XICDRVM0/XICDRV0/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV0/XISW0/XIN1/MM0 VREF<2> ZP<1> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV0/XISW0/XIN0/MM0 VREF<2> ZP<1> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV0/XISW1/XIN1/MM0 VREF<1> ZMID<1> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV0/XISW1/XIN0/MM0 VREF<1> ZMID<1> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV0/XISW2/XIN1/MM0 VREF<0> ZM<1> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV0/XISW2/XIN0/MM0 VREF<0> ZM<1> VOR<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV2/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV2/XITIE0/net5 XISAR0/XIAFE0/XICDRVM0/XICDRV2/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV2/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV2/XITIE0/net6 XISAR0/XIAFE0/XICDRVM0/XICDRV2/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV2/XISW0/XIN1/MM0 VREF<2> ZP<3> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV2/XISW0/XIN0/MM0 VREF<2> ZP<3> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV2/XISW1/XIN1/MM0 VREF<1> ZMID<3> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV2/XISW1/XIN0/MM0 VREF<1> ZMID<3> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV2/XISW2/XIN1/MM0 VREF<0> ZM<3> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV2/XISW2/XIN0/MM0 VREF<0> ZM<3> VOR<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV1/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV1/XITIE0/net5 XISAR0/XIAFE0/XICDRVM0/XICDRV1/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV1/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV1/XITIE0/net6 XISAR0/XIAFE0/XICDRVM0/XICDRV1/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV1/XISW0/XIN1/MM0 VREF<2> ZP<2> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV1/XISW0/XIN0/MM0 VREF<2> ZP<2> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV1/XISW1/XIN1/MM0 VREF<1> ZMID<2> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV1/XISW1/XIN0/MM0 VREF<1> ZMID<2> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV1/XISW2/XIN1/MM0 VREF<0> ZM<2> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV1/XISW2/XIN0/MM0 VREF<0> ZM<2> VOR<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV4/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV4/XITIE0/net5 XISAR0/XIAFE0/XICDRVM0/XICDRV4/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV4/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV4/XITIE0/net6 XISAR0/XIAFE0/XICDRVM0/XICDRV4/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV4/XISW0/XIN1/MM0 VREF<2> ZP<5> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV4/XISW0/XIN0/MM0 VREF<2> ZP<5> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV4/XISW1/XIN1/MM0 VREF<1> ZMID<5> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV4/XISW1/XIN0/MM0 VREF<1> ZMID<5> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV4/XISW2/XIN1/MM0 VREF<0> ZM<5> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV4/XISW2/XIN0/MM0 VREF<0> ZM<5> VOR<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV5/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV5/XITIE0/net5 XISAR0/XIAFE0/XICDRVM0/XICDRV5/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV5/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV5/XITIE0/net6 XISAR0/XIAFE0/XICDRVM0/XICDRV5/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV5/XISW0/XIN1/MM0 VREF<2> ZP<6> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV5/XISW0/XIN0/MM0 VREF<2> ZP<6> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV5/XISW1/XIN1/MM0 VREF<1> ZMID<6> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV5/XISW1/XIN0/MM0 VREF<1> ZMID<6> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV5/XISW2/XIN1/MM0 VREF<0> ZM<6> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV5/XISW2/XIN0/MM0 VREF<0> ZM<6> VOR<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV6/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV6/XITIE0/net5 XISAR0/XIAFE0/XICDRVM0/XICDRV6/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV6/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV6/XITIE0/net6 XISAR0/XIAFE0/XICDRVM0/XICDRV6/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV6/XISW0/XIN1/MM0 VREF<2> ZP<7> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVM0/XICDRV6/XISW0/XIN0/MM0 VREF<2> ZP<7> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVM0/XICDRV6/XISW1/XIN1/MM0 VREF<1> ZMID<7> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVM0/XICDRV6/XISW1/XIN0/MM0 VREF<1> ZMID<7> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVM0/XICDRV6/XISW2/XIN1/MM0 VREF<0> ZM<7> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVM0/XICDRV6/XISW2/XIN0/MM0 VREF<0> ZM<7> VOR<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVM0/XICDRV7/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV7/XITIE0/net5 XISAR0/XIAFE0/XICDRVM0/XICDRV7/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV7/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVM0/XICDRV7/XITIE0/net6 XISAR0/XIAFE0/XICDRVM0/XICDRV7/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVM0/XICDRV7/XISW0/XIN1/MM0 VREF<2> ZP<8> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVM0/XICDRV7/XISW0/XIN0/MM0 VREF<2> ZP<8> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVM0/XICDRV7/XISW1/XIN1/MM0 VREF<1> ZMID<8> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVM0/XICDRV7/XISW1/XIN0/MM0 VREF<1> ZMID<8> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVM0/XICDRV7/XISW2/XIN1/MM0 VREF<0> ZM<8> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVM0/XICDRV7/XISW2/XIN0/MM0 VREF<0> ZM<8> VOR<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVP0/XICDRV3/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV3/XITIE0/net5 XISAR0/XIAFE0/XICDRVP0/XICDRV3/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV3/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV3/XITIE0/net6 XISAR0/XIAFE0/XICDRVP0/XICDRV3/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV3/XISW0/XIN1/MM0 VREF<2> ZM<4> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV3/XISW0/XIN0/MM0 VREF<2> ZM<4> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV3/XISW1/XIN1/MM0 VREF<1> ZMID<4> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV3/XISW1/XIN0/MM0 VREF<1> ZMID<4> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV3/XISW2/XIN1/MM0 VREF<0> ZP<4> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV3/XISW2/XIN0/MM0 VREF<0> ZP<4> VOL<3> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV0/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV0/XITIE0/net5 XISAR0/XIAFE0/XICDRVP0/XICDRV0/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV0/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV0/XITIE0/net6 XISAR0/XIAFE0/XICDRVP0/XICDRV0/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV0/XISW0/XIN1/MM0 VREF<2> ZM<1> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV0/XISW0/XIN0/MM0 VREF<2> ZM<1> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV0/XISW1/XIN1/MM0 VREF<1> ZMID<1> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV0/XISW1/XIN0/MM0 VREF<1> ZMID<1> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV0/XISW2/XIN1/MM0 VREF<0> ZP<1> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV0/XISW2/XIN0/MM0 VREF<0> ZP<1> VOL<0> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV2/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV2/XITIE0/net5 XISAR0/XIAFE0/XICDRVP0/XICDRV2/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV2/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV2/XITIE0/net6 XISAR0/XIAFE0/XICDRVP0/XICDRV2/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV2/XISW0/XIN1/MM0 VREF<2> ZM<3> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV2/XISW0/XIN0/MM0 VREF<2> ZM<3> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV2/XISW1/XIN1/MM0 VREF<1> ZMID<3> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV2/XISW1/XIN0/MM0 VREF<1> ZMID<3> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV2/XISW2/XIN1/MM0 VREF<0> ZP<3> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV2/XISW2/XIN0/MM0 VREF<0> ZP<3> VOL<2> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV1/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV1/XITIE0/net5 XISAR0/XIAFE0/XICDRVP0/XICDRV1/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV1/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV1/XITIE0/net6 XISAR0/XIAFE0/XICDRVP0/XICDRV1/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV1/XISW0/XIN1/MM0 VREF<2> ZM<2> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV1/XISW0/XIN0/MM0 VREF<2> ZM<2> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV1/XISW1/XIN1/MM0 VREF<1> ZMID<2> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV1/XISW1/XIN0/MM0 VREF<1> ZMID<2> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV1/XISW2/XIN1/MM0 VREF<0> ZP<2> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV1/XISW2/XIN0/MM0 VREF<0> ZP<2> VOL<1> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV4/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV4/XITIE0/net5 XISAR0/XIAFE0/XICDRVP0/XICDRV4/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV4/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV4/XITIE0/net6 XISAR0/XIAFE0/XICDRVP0/XICDRV4/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV4/XISW0/XIN1/MM0 VREF<2> ZM<5> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV4/XISW0/XIN0/MM0 VREF<2> ZM<5> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV4/XISW1/XIN1/MM0 VREF<1> ZMID<5> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV4/XISW1/XIN0/MM0 VREF<1> ZMID<5> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV4/XISW2/XIN1/MM0 VREF<0> ZP<5> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV4/XISW2/XIN0/MM0 VREF<0> ZP<5> VOL<4> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV5/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV5/XITIE0/net5 XISAR0/XIAFE0/XICDRVP0/XICDRV5/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV5/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV5/XITIE0/net6 XISAR0/XIAFE0/XICDRVP0/XICDRV5/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV5/XISW0/XIN1/MM0 VREF<2> ZM<6> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV5/XISW0/XIN0/MM0 VREF<2> ZM<6> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV5/XISW1/XIN1/MM0 VREF<1> ZMID<6> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV5/XISW1/XIN0/MM0 VREF<1> ZMID<6> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV5/XISW2/XIN1/MM0 VREF<0> ZP<6> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV5/XISW2/XIN0/MM0 VREF<0> ZP<6> VOL<5> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV6/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV6/XITIE0/net5 XISAR0/XIAFE0/XICDRVP0/XICDRV6/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV6/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV6/XITIE0/net6 XISAR0/XIAFE0/XICDRVP0/XICDRV6/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV6/XISW0/XIN1/MM0 VREF<2> ZM<7> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVP0/XICDRV6/XISW0/XIN0/MM0 VREF<2> ZM<7> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVP0/XICDRV6/XISW1/XIN1/MM0 VREF<1> ZMID<7> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVP0/XICDRV6/XISW1/XIN0/MM0 VREF<1> ZMID<7> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVP0/XICDRV6/XISW2/XIN1/MM0 VREF<0> ZP<7> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVP0/XICDRV6/XISW2/XIN0/MM0 VREF<0> ZP<7> VOL<6> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXISAR0/XIAFE0/XICDRVP0/XICDRV7/XITIE0/XIN1/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV7/XITIE0/net5 XISAR0/XIAFE0/XICDRVP0/XICDRV7/XITIE0/net5 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV7/XITIE0/XIN0/MM0 XISAR0/XIAFE0/XICDRVP0/XICDRV7/XITIE0/net6 XISAR0/XIAFE0/XICDRVP0/XICDRV7/XITIE0/net6 VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=2 
MXISAR0/XIAFE0/XICDRVP0/XICDRV7/XISW0/XIN1/MM0 VREF<2> ZM<8> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVP0/XICDRV7/XISW0/XIN0/MM0 VREF<2> ZM<8> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVP0/XICDRV7/XISW1/XIN1/MM0 VREF<1> ZMID<8> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVP0/XICDRV7/XISW1/XIN0/MM0 VREF<1> ZMID<8> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVP0/XICDRV7/XISW2/XIN1/MM0 VREF<0> ZP<8> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXISAR0/XIAFE0/XICDRVP0/XICDRV7/XISW2/XIN0/MM0 VREF<0> ZP<8> VOL<7> VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
RXISAR0/XIAFE0/XICAPM0/XI7<99>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<98>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<97>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<96>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<95>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<94>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<93>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<92>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<91>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<90>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<89>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<88>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<87>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<86>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<85>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<84>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<83>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<82>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<81>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<80>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<79>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<78>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<77>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<76>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<75>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<74>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<73>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<72>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<71>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<70>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<69>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<68>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<67>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<66>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<65>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<64>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<63>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<62>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<61>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<60>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<59>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<58>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<57>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<56>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<55>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<54>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<53>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<52>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<51>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<50>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<49>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<48>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<47>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<46>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<45>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<44>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<43>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<42>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<41>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<40>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<39>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<38>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<37>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<36>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<35>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<34>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<33>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<32>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<31>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<30>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<29>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<28>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<27>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<26>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<25>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<24>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<23>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<22>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<21>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<20>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<19>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<18>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<17>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<16>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<15>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<14>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<13>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<12>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<11>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<10>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<9>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<8>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<7>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<6>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<5>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<4>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<3>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<2>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<1>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI7<0>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<52>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<51>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<50>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<49>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<48>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<47>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<46>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<45>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<44>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<43>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<42>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<41>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<40>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<39>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<38>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<37>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<36>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<35>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<34>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<33>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<32>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<31>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<30>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<29>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<28>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<27>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<26>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<25>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<24>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<23>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<22>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<21>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<20>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<19>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<18>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<17>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<16>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<15>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<14>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<13>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<12>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<11>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<10>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<9>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<8>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<7>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<6>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<5>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<4>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<3>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<2>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<1>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI6<0>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<27>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<26>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<25>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<24>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<23>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<22>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<21>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<20>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<19>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<18>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<17>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<16>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<15>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<14>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<13>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<12>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<11>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<10>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<9>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<8>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<7>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<6>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<5>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<4>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<3>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<2>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<1>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI5<0>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<15>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<14>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<13>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<12>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<11>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<10>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<9>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<8>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<7>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<6>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<5>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<4>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<3>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<2>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<1>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI4<0>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI3<7>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI3<6>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI3<5>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI3<4>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI3<3>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI3<2>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI3<1>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI3<0>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI2<3>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI2<2>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI2<1>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI2<0>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI1<1>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI1<0>/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XIC0_0/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPM0/XI0/RR0 SAMPM SAMPM RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<99>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<98>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<97>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<96>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<95>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<94>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<93>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<92>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<91>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<90>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<89>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<88>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<87>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<86>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<85>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<84>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<83>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<82>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<81>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<80>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<79>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<78>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<77>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<76>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<75>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<74>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<73>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<72>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<71>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<70>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<69>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<68>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<67>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<66>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<65>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<64>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<63>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<62>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<61>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<60>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<59>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<58>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<57>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<56>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<55>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<54>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<53>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<52>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<51>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<50>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<49>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<48>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<47>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<46>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<45>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<44>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<43>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<42>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<41>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<40>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<39>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<38>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<37>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<36>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<35>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<34>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<33>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<32>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<31>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<30>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<29>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<28>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<27>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<26>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<25>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<24>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<23>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<22>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<21>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<20>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<19>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<18>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<17>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<16>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<15>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<14>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<13>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<12>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<11>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<10>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<9>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<8>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<7>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<6>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<5>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<4>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<3>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<2>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<1>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI7<0>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<52>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<51>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<50>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<49>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<48>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<47>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<46>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<45>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<44>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<43>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<42>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<41>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<40>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<39>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<38>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<37>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<36>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<35>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<34>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<33>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<32>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<31>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<30>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<29>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<28>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<27>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<26>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<25>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<24>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<23>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<22>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<21>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<20>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<19>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<18>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<17>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<16>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<15>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<14>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<13>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<12>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<11>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<10>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<9>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<8>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<7>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<6>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<5>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<4>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<3>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<2>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<1>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI6<0>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<27>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<26>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<25>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<24>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<23>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<22>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<21>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<20>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<19>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<18>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<17>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<16>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<15>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<14>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<13>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<12>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<11>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<10>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<9>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<8>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<7>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<6>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<5>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<4>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<3>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<2>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<1>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI5<0>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<15>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<14>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<13>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<12>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<11>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<10>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<9>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<8>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<7>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<6>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<5>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<4>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<3>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<2>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<1>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI4<0>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI3<7>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI3<6>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI3<5>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI3<4>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI3<3>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI3<2>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI3<1>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI3<0>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI2<3>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI2<2>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI2<1>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI2<0>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI1<1>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI1<0>/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XIC0_0/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
RXISAR0/XIAFE0/XICAPP0/XI0/RR0 SAMPP SAMPP RESM4 r=0.0604 w=3.2e-08 l=3.2e-08 m=1 
MXXSAMP0/XIBUFB0/XIN0/MM0 XXSAMP0/out_int<0> CLKPRB_SAMP VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXXSAMP0/XIBUFB0/XIP0/MM0 XXSAMP0/out_int<0> CLKPRB_SAMP VDDSAMP VDDSAMP P1LVT m=1 l=1.8e-08 nfin=4 nf=8 
MXXSAMP0/XIBUFA0/XIN0/MM0 XXSAMP0/in_int<0> CLK VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=16 
MXXSAMP0/XIBUFA0/XIP0/MM0 XXSAMP0/in_int<0> CLK VDDSAMP VDDSAMP P1LVT m=1 l=1.8e-08 nfin=4 nf=16 
MXXSAMP0/XISWP<3>/XIN1/MM0 INP CLKPRB_SAMP SAMPP VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWP<3>/XIN0/MM0 INP CLKPRB_SAMP SAMPP VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWP<2>/XIN1/MM0 INP CLKPRB_SAMP SAMPP VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWP<2>/XIN0/MM0 INP CLKPRB_SAMP SAMPP VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWP<1>/XIN1/MM0 INP CLKPRB_SAMP SAMPP VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWP<1>/XIN0/MM0 INP CLKPRB_SAMP SAMPP VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWP<0>/XIN1/MM0 INP CLKPRB_SAMP SAMPP VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWP<0>/XIN0/MM0 INP CLKPRB_SAMP SAMPP VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWN<3>/XIN1/MM0 INM CLKPRB_SAMP SAMPM VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWN<3>/XIN0/MM0 INM CLKPRB_SAMP SAMPM VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWN<2>/XIN1/MM0 INM CLKPRB_SAMP SAMPM VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWN<2>/XIN0/MM0 INM CLKPRB_SAMP SAMPM VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWN<1>/XIN1/MM0 INM CLKPRB_SAMP SAMPM VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWN<1>/XIN0/MM0 INM CLKPRB_SAMP SAMPM VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWN<0>/XIN1/MM0 INM CLKPRB_SAMP SAMPM VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XISWN<0>/XIN0/MM0 INM CLKPRB_SAMP SAMPM VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=4 
MXXSAMP0/XIBUFB1/XIN0/MM0 ICLK XXSAMP0/out_int<0> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=32 
MXXSAMP0/XIBUFB1/XIP0/MM0 ICLK XXSAMP0/out_int<0> VDDSAMP VDDSAMP P1LVT m=1 l=1.8e-08 nfin=4 nf=32 
MXXSAMP0/XIBUFA1/XIN0/MM0 CLKPRB_SAMP XXSAMP0/in_int<0> VSS VSS N1LVT m=1 l=1.8e-08 nfin=4 nf=24 
MXXSAMP0/XIBUFA1/XIP0/MM0 CLKPRB_SAMP XXSAMP0/in_int<0> VDDSAMP VDDSAMP P1LVT m=1 l=1.8e-08 nfin=4 nf=24 
.ends


